// VGA Controller
// James Kaden Cassidy 
// kacassidy@hmc.edu
// 11/12/2025

module state_communicator #(
    
    )(

    );

    game_state_pkg::game_state_t current_game_state, next_game_state;
    


endmodule