// Game Encoder
// James Kaden Cassidy 
// kacassidy@hmc.edu
// 11/12/2025

module game_encoder (
    output  logic                               GAME_new_frame_ready, // not driven here
    output  game_state_pkg::game_state_t        GAME_next_frame
);

    import game_state_pkg::*;
       

endmodule
