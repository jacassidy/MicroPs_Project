// VGA Controller
// James Kaden Cassidy 
// kacassidy@hmce.edu
// 11/8/2025