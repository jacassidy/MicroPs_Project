// Parameters
// James Kaden Cassidy 
// kacassidy@hmc.edu
// 11/13/2025

`ifndef PARAMETERS
`define PARAMETERS
    `define DEBUG
    `define COLORS 3

`endif